module ID_tb();
	initial begin
		$display("\n---------------------------");
		$display("Teste de integracao (ID)");
		$display("Total de testes: ");
	end
endmodule