module signal_generator_tb;
endmodule
