module signal_generator(
	input 	wire[2:0]	type,
	input 	wire[4:0]	op,
	output 	reg 		byPass
	);
	//meudeus oq será q vai acontecer aqui gzus
	always @ (*) begin
		
	end
endmodule
