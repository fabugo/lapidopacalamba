module EX();
endmodule
