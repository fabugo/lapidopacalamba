module forward_unit_tb;
endmodule
