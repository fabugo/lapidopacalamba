module WB();

endmodule
