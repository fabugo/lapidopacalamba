module mx_a_tb;
endmodule
