module processor;

    unit_control uc(CLK,
                    type,
                    op);

endmodule
