module IF_ID_tb;
endmodule
