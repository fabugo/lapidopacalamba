module mi_rb_tb();
	//Cria a memória
	//memory_instruction u1();

	initial begin
		$display("\n---------------------------");
		$display("Teste de integracao (MI - RB)");
		$display("Total de testes: ");
	end
endmodule