module ex_tb();
	initial begin
		$display("\n---------------------------");
		$display("Teste de integracao (EX)");
		$display("Total de testes: ");
	end
endmodule