module WB_tb;
endmodule
