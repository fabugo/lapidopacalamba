module reg_EXMEM_WB_tb;
endmodule
