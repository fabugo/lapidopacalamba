module unit_control();
endmodule