module mx_b_tb;
endmodule
