module wb_tb();
	initial begin
		$display("\n---------------------------");
		$display("Teste de integracao (WB)");
		$display("Total de testes: ");
	end
endmodule