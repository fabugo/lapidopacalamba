module EX_MEM_tb;
endmodule
