module memory_instruction(
			input 	wire[31:0]	in,
			input 	wire		W_MI,
			output 	reg[31:0]	out);

	reg[31:0] 	instruction[0:1024];

	always @() begin
	end

endmodule