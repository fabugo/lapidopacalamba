module WB();
endmodule
