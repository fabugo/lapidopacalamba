module reg_IFID_EXMEM_tb;
endmodule
