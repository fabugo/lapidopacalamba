module if_tb();
	initial begin
		$display("\n---------------------------");
		$display("Teste de integracao (IF)");
		$display("Total de testes: ");
	end
endmodule